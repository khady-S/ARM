----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/05/2025 10:10:05 PM
-- Design Name: 
-- Module Name: memoire_instruction - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity memoire_instruction is
    Port (
        A  : in  STD_LOGIC_VECTOR(31 downto 0);
        RD : out STD_LOGIC_VECTOR(31 downto 0)
    );
end memoire_instruction;

architecture Behavioral of memoire_instruction is
    type ramtype is array (0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
    
    --PROGRAMME DE TEST SHIFTED REGISTER
    signal mem : ramtype := (
        0  => "11100000010000000000000000000000",
        1  => "11100010100000000010000000000101",
        2  => "11100010100000000011000000001100",
        3  => "11100010010000110111000000001001",
        4  => "11100001100001110100000000000010",
        5  => "11100000000000110101000000000100",
        6  => "11100000100001010101000000000100",
        7  => "11100000010101011000000000000111",
        8  => "11100000010100111000000000000100",
        9  => "11100010100000000101000000000000",
        10 => "11100000010101111000000000000010",
        11 => "10110010100001010111000000000001",
        12 => "11100000010001110111000000000010",
        13 => "11100101100000110111000001010100",
        14 => "11100101100100000010000001100000",
        15 => "11100000100010000101000000000000",
        16 => "11100010100000000010000000001110",
        17 => "11100010100000000010000000001101",
        18 => "11100010100000000010000000001010",
        19 => "11100101100000000010000001100100",
    
        -- Test 1: LSL (Logical Shift Left)
--        0  => "11100011101000000000000000001000",  -- MOV R0, #8
--        1  => "11100000100000000001000010000000",  -- ADD R1, R0, R0, LSL #1 (8 << 1 = 16, R1 = 8 + 16 = 24)

        
--        -- Test 2: LSL avec shift amount plus grand
--        2  => "11100011101000000010000000000001",  -- MOV R2, #1
--        3  => "11100000010000000011001000100010",  -- ADD R3, R0, R2, LSL #4 (1 << 4 = 16, R3 = 8 + 16 = 24)
        
--        -- Test 3: LSR (Logical Shift Right)
--        4  => "11100011101000000100000010000000",  -- MOV R4, #128 (0x80)
--        5  => "11100000010000000101001000100100",  -- ADD R5, R0, R4, LSR #4 (128 >> 4 = 8, R5 = 8 + 8 = 16)
        
--        -- Test 4: ASR (Arithmetic Shift Right) avec nombre n�gatif
--        6  => "11100011111000000110111111111111",  -- MVN R6, #0 (R6 = -1 = 0xFFFFFFFF)
--        7  => "11100000010000000111001101000110",  -- ADD R7, R0, R6, ASR #2 (-1 >> 2 = -1, R7 = 8 + (-1) = 7)
        
--        -- Test 5: ROR (Rotate Right)
--        8  => "11100011101000001000000010000000",  -- MOV R8, #128
--        9  => "11100000010000001001010000110000", -- ADD R9, R0, R8, ROR #1 (rotate 128 = 64, R9 = 8 + 64 = 72)
        
--        -- Test 6: Sans shift (v�rifier que �a marche toujours)
--        10 => "11100011101000001010000000000101",  -- MOV R10, #5
--        11 => "11100000010010101011000000001010",  -- ADD R11, R10, R10 (5 + 5 = 10)
        
--  -- =====================================================================
--        -- SECTION 2: TESTS CMP (Compare)
--        -- =====================================================================
        
--        -- Test 7: CMP �galit� (R12 = R13) -> Z=1, C=1
--        12 => "11100011101000001100000000001010",  -- MOV R12, #10
--        13 => "11100011101000001101000000001010",  -- MOV R13, #10
--        14 => "11100001010111000000000000001101",  -- CMP R12, R13 (10-10=0, Z=1, C=1)
        
--        -- Test 8: CMP plus petit (5 < 15) -> N=1, C=0
--        15 => "11100011101000001110000000000101",  -- MOV R14, #5
--        16 => "11100011101000000000000000001111",  -- MOV R0, #15 (r�utilise R0)
--        17 => "11100001010111100000000000000000",  -- CMP R14, R0 (5-15=-10, N=1, C=0)
        
--        -- Test 9: CMP plus grand (20 > 3) -> C=1, N=0, Z=0
--        18 => "11100011101000000001000000010100",  -- MOV R1, #20
--        19 => "11100011101000000010000000000011",  -- MOV R2, #3
--        20 => "11100001010100010000000000000010",  -- CMP R1, R2 (20-3=17, C=1)
        
--        -- Test 10: CMP avec z�ro (0 = 0) -> Z=1, C=1
--        21 => "11100011101000000011000000000000",  -- MOV R3, #0
--        22 => "11100011101000000100000000000000",  -- MOV R4, #0
--        23 => "11100001010100110000000000000100",  -- CMP R3, R4 (0-0=0, Z=1, C=1)
        
--        -- Test 11: V�rifier que CMP ne modifie pas les registres
--        24 => "11100011101000000101000000100000",  -- MOV R5, #32
--        25 => "11100011101000000110000000010000",  -- MOV R6, #16
--        26 => "11100001010101010000000000000110",  -- CMP R5, R6 (32-16=16, pas d'�criture)
----        27 => "11100000010001010111000000000110",  -- ADD R7, R5, R6 (V�rif: R5=32, R6=16 -> R7=48)
        
--        -- Test 12: CMP avec nombre n�gatif
--        30 => "11100011111000001000000000001010",  -- MVN R8, #10 (R8 = -11 = 0xFFFFFFF5)
--        31 => "11100011101000001001000000000101",  -- MOV R9, #5
--        32 => "11100001010110000000000000001001",  -- CMP R8, R9 (n�gatif < positif, N=1)
        
        others => (others => '0')
    );
    
begin
    RD <= mem(to_integer(unsigned(A(6 downto 2))));
end Behavioral;

---

