----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10/09/2025 11:33:37 AM
-- Design Name: 
-- Module Name: Data_Memory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Data_Memory is
    Port (
        -- Entr�es
        CLK : in STD_LOGIC;                       -- Signal d'horloge
        MemWrite : in STD_LOGIC;                  -- Activation �criture (1 = �crire)
        A : in STD_LOGIC_VECTOR(31 downto 0);     -- Adresse m�moire
        WD : in STD_LOGIC_VECTOR(31 downto 0);    -- Donn�e � �crire
        
        -- Sortie
        RD : out STD_LOGIC_VECTOR(31 downto 0)    -- Donn�e lue
    );
end Data_Memory;

architecture Behavioral of Data_Memory is
    -- D�claration de la m�moire : 64 cases de 32 bits
    type ramtype is array (0 to 63) of STD_LOGIC_VECTOR(31 downto 0);
    signal mem : ramtype := (others => (others => '0'));  -- Initialisation � z�ro
    
begin

    -- Processus d'�criture synchrone
    process(CLK) 
    begin
        -- Sur front montant d'horloge
        if rising_edge(CLK) then
            -- Si �criture activ�e
            if MemWrite = '1' then 
            -- �crire WD � l'adresse A (seuls 6 bits utilis�s)
                mem(to_integer(unsigned(A(5 downto 0)))) <= WD;
            end if;
        end if;
    end process;

    -- Processus de lecture asynchrone

        -- Lire toujours la donn�e � l'adresse A
        RD <= mem(to_integer(unsigned(A(5 downto 0))));

end Behavioral;